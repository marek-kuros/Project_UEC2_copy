module char_rom_16x16(
    input  logic [7:0] char_xy,
    input  logic [3:0] char_line,
    output logic [10:0] char_code
);

typedef bit [7:0] array_byte;

logic [3:0] x_pos;
logic [3:0] y_pos;

array_byte [15:0][15:0] array_of_letters = '{
                        '{"T", "R", "Y", "B", " ", " ", " ", "G", "R", "Y", "", "", "", "", "", ""},
                        '{"", "", "", "", "", "", "", "", "", "", "", "", "", "", "", ""},
                        '{"", "", "", "", "", "", "", "", "", "", "", "", "", "", "", ""},
                        '{"", "", "", "", "", "", "", "", "", "", "", "", "", "", "", ""},
                        '{"", "", "", "", "", "", "", "", "", "", "", "", "", "", "", ""},
                        '{"", "", "", "", "", "", "", "", "", "", "", "", "", "", "", ""},
                        '{"", "", "", "", "", "", "", "", "", "", "", "", "", "", "", ""},
                        '{"S", "I", "N", "G", "L", "E", "", "", "", "", "", "", "", "", "", ""},
                        '{"", "", "", "", "", "", "", "", "", "", "", "", "", "", "", ""},
                        '{"", "", "", "", "", "", "", "", "", "", "", "", "", "", "", ""},
                        '{"", "", "", "", "", "", "", "", "", "", "", "", "", "", "", ""},
                        '{"", "", "", "", "", "", "", "", "", "", "", "", "", "", "", ""},
                        '{"", "", "", "", "", "", "", "", "", "", "", "", "", "", "", ""},
                        '{"", "", "", "", "", "", "", "", "", "", "", "", "", "", "", ""},
                        '{"M", "U", "L", "T", "I", "", "", "", "", "", "", "", "", "", "", ""},
                        '{"", "", "", "", "", "", "", "", "", "", "", "", "", "", "", ""}
                    };
always_comb begin
    x_pos = char_xy[7:4];
    y_pos = char_xy[3:0];
end

logic [10:4] value;

always_comb begin
    value = array_of_letters[15 - x_pos][15 - y_pos];
    char_code[10:0] = {value, char_line};
end

endmodule